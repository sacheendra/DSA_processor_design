module alu_mov(A, B, Y);

input [31:0] A, B;
output [31:0] Y;

assign Y = B;
endmodule