module fetch(
    input clk,
    input [31:0] br_pc,
    input Br,
    input [31:0] pc_pred,
    output reg [31:0] instr
    );
    
    reg [31:0] pc = 31'd0;
    
    reg [31:0] mem [10:0];
    wire pred = 1'b0;

    initial begin
        mem[32'd0] = 32'b01001001000100000000000000000001; //sub
        mem[32'd1] = 32'b01011101000100000000000000000001; //cmp
        mem[32'd2] = 32'b00100100000000000000000000000000; //branch
        mem[32'd3] = 32'b00000110000100000000000000000011; //add
		  mem[32'd4] = 32'b00111001001100001000010000000010; //ldr
		  mem[32'd5] = 32'b00000110000000010000000000000011; //add
    end
    
    always @(posedge clk) begin
        instr <= mem[pc];
    end
    
    always @(negedge clk) begin
	if(instr[29] == 1 && instr[28] == 0) begin
		pred = 1'b1;
	end
	case({Br, pred})
	2'b00: pc <= pc+32'd1;
	2'b01: pc <= br_pc;
	2'b10: pc <= pc_pred;
	2'b11: pc <= br_pc;
        if(Br) begin
	pc <= br_pc;
	end
	else begin
	pc <= pc+32'd1;
	end
    end

endmodule

mem[32'd0] = 32'b10111001101100000000000000001010;//32'b01001001000100000000000000000001; //sub
        mem[32'd1] = 32'b10111001110000000000000000010100; //cmp
		  mem[32'd2] = 32'd0;
		  mem[32'd3] = 32'd0;
        mem[32'd4] = 32'b00011100110000000000000000001100; //branch
        mem[32'd5] = 32'b11000110110111010000000000000010; //add
		  mem[32'd6] = 32'b00100101000000000000000000000100; //ldr
		  mem[32'd7] = 32'b00100100000000000000000000001011; //add
		  mem[32'd8] = 32'b01001110110011100000000000001011;
		  mem[32'd9] = 32'd0;
		  mem[32'd10] = 32'd0;
		  mem[32'd11] = 32'b11001010111011100000000000000111;
		  mem[32'd12] = 32'b00110010000000000000000000000100;
		  mem[32'd13] = 32'b00000110111011110000000000001101;
		  mem[32'd14] = 32'd0;
		  mem[32'd15] = 32'd0; 
		  mem[32'd16] = 32'd0;
		  mem[32'd17] = 32'd0;
		  mem[32'd18] = 32'd0;